`include "../include/define.svh"


module top (
    input clk,
    input rst,
    
);
    
endmodule